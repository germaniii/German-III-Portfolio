//GERMAN E FELISARTA III 16101002	CpE 3101L

module hexaDigit(Hex, DP, SSeg);
	
	input wire [3:0]Hex;
	input wire DP;
	output reg [7:0]SSeg;
	
	always @ (*)
		begin
				case ({DP, Hex})
					5'b00000 : SSeg = 8'b0111111;
					5'b00001 : SSeg = 8'b0000110;
					5'b00010 : SSeg = 8'b1011011;
					5'b00011 : SSeg = 8'b1001111;
					5'b00100 : SSeg = 8'b1100110;
					5'b00101 : SSeg = 8'b1101101;
					5'b00110 : SSeg = 8'b1111101;
					5'b00111 : SSeg = 8'b0000111;
					5'b01000 : SSeg = 8'b1111111;
					5'b01001 : SSeg = 8'b1101111;
					5'b01010 : SSeg = 8'b1110111;
					5'b01011 : SSeg = 8'b1111100;
					5'b01100 : SSeg = 8'b0111001;
					5'b01101 : SSeg = 8'b1011110;
					5'b01110 : SSeg = 8'b1111001;
					5'b01111 : SSeg = 8'b1110001;
					default : SSeg = 8'b0000000;
					
				endcase
		end
		
endmodule

				
/*				  GFEDCBA
		0000 - 0 - 0111111
		0001 - 1 - 0000110
		0010 - 2 - 1011011
		0011 - 3 - 1001111
		0100 - 4 - 1100110
		0101 - 5 - 1101101
		0110 - 6 - 1111101
		0111 - 7 - 0000111
		1000 - 8 - 1111111
		1001 - 9 - 1101111
		1010 - A - 1110111
		1011 - B - 1111100
		1100 - C - 0111001
		1101 - D - 1011110
		1110 - E - 1111001
		1111 - F - 1110001
	*/